library verilog;
use verilog.vl_types.all;
entity FIFO_tb is
end FIFO_tb;
